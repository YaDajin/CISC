LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY MUX3_1 IS
PORT(
	INBUS,RAMOUT,FEN2OUT:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	SW_B,RAM_B:IN STD_LOGIC;
	DBUS:OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END MUX3_1;

ARCHITECTURE A OF MUX3_1 IS
BEGIN
    PROCESS
     BEGIN 
       IF(SW_B='0') THEN     			
            DBUS<=INBUS;
	   ELSIF(RAM_B='0')THEN 
			DBUS<=RAMOUT;			
	   ELSE
			DBUS<=FEN2OUT;
		END IF;
    END PROCESS;
END A;

