LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY ROM IS 
PORT(
	DOUT:OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	ADDR:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	CS_I:IN STD_LOGIC
);
END ROM;
ARCHITECTURE A OF ROM IS

--  ע�Ƿ���    ָ���ʽ(OP)    Rs Rd     addr   
--    MOV            0001       XX Rd    XXXXXXXX
--    INT            0010       XX Rd    XXXXXXXX
--    TEST           0011       Rs XX    XXXXXXXX
--    JB             0100       XX XX     addr
--    MUL            0101       Rs Rd    XXXXXXXX
--    ADD            0110       Rs Rd    XXXXXXXX
--    DEC            0111       XX Rd    XXXXXXXX
--    JZ             1000       XX XX     addr
--    OUT            1001       Rs XX    XXXXXXXX
--    JMP            1010       XX XX     addr
BEGIN
	DOUT<="0001001100000000" WHEN ADDR=x"00" AND CS_I='0' ELSE--MOV R3,0H
          "0001000100000101" WHEN ADDR=x"01" AND CS_I='0' ELSE--MOV R1,5H
          "0011010000000000" WHEN ADDR=x"02" AND CS_I='0' ELSE--L1:TEST R1
		  "1000000000001011" WHEN ADDR=x"03" AND CS_I='0' ELSE--JZ L2
          "0010001000000000" WHEN ADDR=x"04" AND CS_I='0' ELSE--INT R2
          "0011100000000000" WHEN ADDR=x"05" AND CS_I='0' ELSE--TEST R2
          "0100000000000010" WHEN ADDR=x"06" AND CS_I='0' ELSE--JB L1
          "0101101000000000" WHEN ADDR=x"07" AND CS_I='0' ELSE--MUL R2,R2
          "0110101100000000" WHEN ADDR=x"08" AND CS_I='0' ELSE--ADD R2,R3
          "0111000100000000" WHEN ADDR=x"09" AND CS_I='0' ELSE--DEC R1
		  "1010000000000010" WHEN ADDR=x"0A" AND CS_I='0' ELSE--JMP L1
		  "1001110000000000" WHEN ADDR=x"0B" AND CS_I='0' ELSE--L2:OUT R3
		  "1010000000001011" WHEN ADDR=x"0C" AND CS_I='0' ELSE--JMP L2
		  "0000000000000000";
END A;

